interface i2c_if(
  inout sda,
  inout scl
);

endinterface
