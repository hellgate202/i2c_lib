interface i2c_int_if(
  input        sda_i,
  output logic sda_o,
  output logic sda_oe,
  input        scl_i,
  output logic scl_o,
  output logic scl_oe
);

endinterface
