package i2c_slave_pkg;

parameter bit [1 : 0] NOP   = 2'b00;
parameter bit [1 : 0] WRITE = 2'b01;
parameter bit [1 : 0] READ  = 2'b10;

endpackage
